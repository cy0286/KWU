module ASR65(d_in,shamt,d_out); //65-bits Arithmetic Shift Right
	input  [64:0] d_in;
	input  [1:0] shamt;
	output [64:0] d_out;
	
	//load mx4 & struct ASR8
	mx4 U0_mx4(d_out[64], d_in[64], d_in[64], d_in[64], d_in[64], shamt);
	mx4 U1_mx4(d_out[63], d_in[63], d_in[64], d_in[64], d_in[64], shamt);
	mx4 U2_mx4(d_out[62], d_in[62], d_in[63], d_in[64], d_in[64], shamt);
	mx4 U3_mx4(d_out[61], d_in[61], d_in[62], d_in[63], d_in[64], shamt);
	mx4 U4_mx4(d_out[60], d_in[60], d_in[61], d_in[62], d_in[63], shamt);
	mx4 U5_mx4(d_out[59], d_in[59], d_in[60], d_in[61], d_in[62], shamt);
	mx4 U6_mx4(d_out[58], d_in[58], d_in[59], d_in[60], d_in[61], shamt);
	mx4 U7_mx4(d_out[57], d_in[57], d_in[58], d_in[59], d_in[60], shamt);
	mx4 U8_mx4(d_out[56], d_in[56], d_in[57], d_in[58], d_in[59], shamt);
	mx4 U9_mx4(d_out[55], d_in[55], d_in[56], d_in[57], d_in[58], shamt);
	mx4 U10_mx4(d_out[54], d_in[54], d_in[55], d_in[56], d_in[57], shamt);
	mx4 U11_mx4(d_out[53], d_in[53], d_in[54], d_in[55], d_in[56], shamt);
	mx4 U12_mx4(d_out[52], d_in[52], d_in[53], d_in[54], d_in[55], shamt);
	mx4 U13_mx4(d_out[51], d_in[51], d_in[52], d_in[53], d_in[54], shamt);
	mx4 U14_mx4(d_out[50], d_in[50], d_in[51], d_in[52], d_in[53], shamt);
	mx4 U15_mx4(d_out[49], d_in[49], d_in[50], d_in[51], d_in[52], shamt);
	mx4 U16_mx4(d_out[48], d_in[48], d_in[49], d_in[50], d_in[51], shamt);
	mx4 U17_mx4(d_out[47], d_in[47], d_in[48], d_in[49], d_in[50], shamt);
	mx4 U18_mx4(d_out[46], d_in[46], d_in[47], d_in[48], d_in[49], shamt);
	mx4 U19_mx4(d_out[45], d_in[45], d_in[46], d_in[47], d_in[48], shamt);
	mx4 U20_mx4(d_out[44], d_in[44], d_in[45], d_in[46], d_in[47], shamt);
	mx4 U21_mx4(d_out[43], d_in[43], d_in[44], d_in[45], d_in[46], shamt);
	mx4 U22_mx4(d_out[42], d_in[42], d_in[43], d_in[44], d_in[45], shamt);
	mx4 U23_mx4(d_out[41], d_in[41], d_in[42], d_in[43], d_in[44], shamt);
	mx4 U24_mx4(d_out[40], d_in[40], d_in[41], d_in[42], d_in[43], shamt);
	mx4 U25_mx4(d_out[39], d_in[39], d_in[40], d_in[41], d_in[42], shamt);
	mx4 U26_mx4(d_out[38], d_in[38], d_in[39], d_in[40], d_in[41], shamt);
	mx4 U27_mx4(d_out[37], d_in[37], d_in[38], d_in[39], d_in[40], shamt);
	mx4 U28_mx4(d_out[36], d_in[36], d_in[37], d_in[38], d_in[39], shamt);
	mx4 U29_mx4(d_out[35], d_in[35], d_in[36], d_in[37], d_in[38], shamt);
	mx4 U30_mx4(d_out[34], d_in[34], d_in[35], d_in[36], d_in[37], shamt);
	mx4 U31_mx4(d_out[33], d_in[33], d_in[34], d_in[35], d_in[36], shamt);
	mx4 U32_mx4(d_out[32], d_in[32], d_in[33], d_in[34], d_in[35], shamt);
	mx4 U33_mx4(d_out[31], d_in[31], d_in[32], d_in[33], d_in[34], shamt);
	mx4 U34_mx4(d_out[30], d_in[30], d_in[31], d_in[32], d_in[33], shamt);
	mx4 U35_mx4(d_out[29], d_in[29], d_in[30], d_in[31], d_in[32], shamt);
	mx4 U36_mx4(d_out[28], d_in[28], d_in[29], d_in[30], d_in[31], shamt);
	mx4 U37_mx4(d_out[27], d_in[27], d_in[28], d_in[29], d_in[30], shamt);
	mx4 U38_mx4(d_out[26], d_in[26], d_in[27], d_in[28], d_in[29], shamt);
	mx4 U39_mx4(d_out[25], d_in[25], d_in[26], d_in[27], d_in[28], shamt);
	mx4 U40_mx4(d_out[24], d_in[24], d_in[25], d_in[26], d_in[27], shamt);
	mx4 U41_mx4(d_out[23], d_in[23], d_in[24], d_in[25], d_in[26], shamt);
	mx4 U42_mx4(d_out[22], d_in[22], d_in[23], d_in[24], d_in[25], shamt);
	mx4 U43_mx4(d_out[21], d_in[21], d_in[22], d_in[23], d_in[24], shamt);
	mx4 U44_mx4(d_out[20], d_in[20], d_in[21], d_in[22], d_in[23], shamt);
	mx4 U45_mx4(d_out[19], d_in[19], d_in[20], d_in[21], d_in[22], shamt);
	mx4 U46_mx4(d_out[18], d_in[18], d_in[19], d_in[20], d_in[21], shamt);
	mx4 U47_mx4(d_out[17], d_in[17], d_in[18], d_in[19], d_in[20], shamt);
	mx4 U48_mx4(d_out[16], d_in[16], d_in[17], d_in[18], d_in[19], shamt);
	mx4 U49_mx4(d_out[15], d_in[15], d_in[16], d_in[17], d_in[18], shamt);
	mx4 U50_mx4(d_out[14], d_in[14], d_in[15], d_in[16], d_in[17], shamt);
	mx4 U51_mx4(d_out[13], d_in[13], d_in[14], d_in[15], d_in[16], shamt);
	mx4 U52_mx4(d_out[12], d_in[12], d_in[13], d_in[14], d_in[15], shamt);
	mx4 U53_mx4(d_out[11], d_in[11], d_in[12], d_in[13], d_in[14], shamt);
	mx4 U54_mx4(d_out[10], d_in[10], d_in[11], d_in[12], d_in[13], shamt);
	mx4 U55_mx4(d_out[9], d_in[9], d_in[10], d_in[11], d_in[12], shamt);
	mx4 U56_mx4(d_out[8], d_in[8], d_in[9], d_in[10], d_in[11], shamt);
	mx4 U57_mx4(d_out[7], d_in[7], d_in[8], d_in[9], d_in[10], shamt);
	mx4 U58_mx4(d_out[6], d_in[6], d_in[7], d_in[8], d_in[9], shamt);
	mx4 U59_mx4(d_out[5], d_in[5], d_in[6], d_in[7], d_in[8], shamt);
	mx4 U60_mx4(d_out[4], d_in[4], d_in[5], d_in[6], d_in[7], shamt);
	mx4 U61_mx4(d_out[3], d_in[3], d_in[4], d_in[5], d_in[6], shamt);
	mx4 U62_mx4(d_out[2], d_in[2], d_in[3], d_in[4], d_in[5], shamt);
	mx4 U63_mx4(d_out[1], d_in[1], d_in[2], d_in[3], d_in[4], shamt);
	mx4 U64_mx4(d_out[0], d_in[0], d_in[1], d_in[2], d_in[3], shamt);
endmodule 